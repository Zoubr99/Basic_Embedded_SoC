//WIP..........